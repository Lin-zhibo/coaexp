`include "ctrl_encode_def.v"

module NPC( PC, NPCOp, IMM, aluout, NPC );  // next pc module
   input  [31:0] PC;        // pc
   input  [2:0]  NPCOp;     // next pc operation
   input  [31:0] IMM;       // immediate
   input  [31:0] aluout;    // alu output
   output reg [31:0] NPC;   // next pc
   
   // default pc += 4
   wire [31:0] PCPLUS4;
   assign PCPLUS4 = PC + 4; // pc + 4
   
   always @(*) begin
      case (NPCOp)
          `NPC_PLUS4:  NPC = PCPLUS4;   // NPC computes addr
          `NPC_BRANCH: NPC = PC+IMM;    //B type, NPC computes addr
          `NPC_JUMP:   NPC = PC+IMM;    //J type, NPC computes 
          `NPC_JALR:   NPC = aluout;
          default:     NPC = PCPLUS4;
      endcase
   end 
   
endmodule
